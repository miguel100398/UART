module UART
module UART_tx
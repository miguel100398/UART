module UART_tx;

endmodule: UART_tx
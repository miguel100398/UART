interface UART_regs_if;

endinterface: UART_regs_if
module UART_tb;

endmodule: UART_tb
module UART_rx;

endmodule: UART_rx
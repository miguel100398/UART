module UART_rx
module UART;

endmodule: UART
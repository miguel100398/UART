
module UART_csr(

);

endmodule: UART_csr
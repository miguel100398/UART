module UART_tb;